module vredis
